-------------------------------------------------------------------------
-- package with basic types
-------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

package p_MR2 is

	subtype reg32 is std_logic_vector(31 downto 0);
	subtype reg16 is std_logic_vector(15 downto 0);
	-- inst_type defines the instructions decodeable by the control unit
	type inst_type is
	(
		ADDU, SUBU, AAND, OOR, XXOR, SSLL, SSRL, ADDIU, ANDI, ORI,
		XORI, LUI, LBU, LW, SB, SW, SLT, SLTU, SLTI, SLTIU, BEQ,
		BGEZ, BLEZ, BNE, J, JALR, JR, RFE, ERET, invalid_instruction
	);

	type microinstruction is record
		CY1: std_logic;	-- command of the first stage
		CY2: std_logic;	--	"	of the second stage
		wula: std_logic;	--	"	of the third stage
		wmdr: std_logic;	--	"	of the fourth stage
		wpc: std_logic;	-- PC write enable
		wreg: std_logic;	-- register bank write enable
		ceRW: std_logic;	-- Chip enable and R_W controls
		rw: std_logic;
		bw: std_logic;	-- Byte-word control (mem write only)
		i: inst_type;	-- operation specification
	end record;

end p_MR2;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- Generic register
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
library IEEE;
use IEEE.std_logic_1164.all;

entity regnbit is
	generic
	(
		N: integer := 16;
		INIT_VALUE: std_logic_vector(31 downto 0) := (others => '0')
	);
	port
	(
		ck, rst, ce: in std_logic;
		D: in std_logic_vector(N-1 downto 0);
		Q: out std_logic_vector(N-1 downto 0)
	);
end regnbit;

architecture regn of regnbit is
begin

	process(ck, rst)
	begin
		if rst = '1' then
			Q <= INIT_VALUE(N-1 downto 0);
		elsif ck'event and ck = '0' then
			if ce = '1' then
				Q <= D;
			end if;
		end if;
	end process;

end regn;

-------------------------------------------------------------------------
-- Register Bank (R0..R31) - 31 GENERAL PURPOSE 16-bit REGISTERS
-------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_UNSIGNED.all;
use work.p_MR2.all;

entity reg_bank is
	port
	(
		ck, rst, wreg: in std_logic;
		AdRs, AdRt, adRD: in std_logic_vector(4 downto 0);
		RD: in reg32;
		R1, R2: out reg32
	);
end reg_bank;

architecture reg_bank of reg_bank is
	type bank is array(0 to 31) of reg32;
	signal reg: bank;
	signal wen: reg32;
begin

	l1: for i in 0 to 31 generate
		wen(i) <= '1' when i/=0 and adRD=i and wreg='1' else '0';
		-- Remember register $0 is the constant 0, not a register.
		-- This is implemented by never enabling writes to register $0
	end generate l1;
	l2: for i in 0 to 28 generate
		rx: entity work.regnbit generic map(N => 32) port map(ck => ck, rst => rst, ce => wen(i), D => RD, Q => reg(i));
	end generate l2;
	--
	--  Beware! Some registers have specific start values - dependent
	-- on code generation. This version is adapted to work with code
	-- generated by the SPIM simulator
	--
	-- SP ---  x10010000 + x800 -- top of stack
	r29: entity work.regnbit generic map(N => 32, INIT_VALUE => x"10010800") port map(ck => ck, rst => rst, ce => wen(29), D => RD, Q => reg(29));
	r30: entity work.regnbit generic map(N => 32) port map(ck => ck, rst => rst, ce => wen(30), D => RD, Q => reg(30));
	-- $ra --
	r31: entity work.regnbit generic map(N => 32) port map(ck => ck, rst => rst, ce => wen(31), D => RD, Q => reg(31));
	R1 <= reg(CONV_INTEGER(AdRs));	-- source1 selection
	R2 <= reg(CONV_INTEGER(AdRt));	-- source2 selection

end reg_bank;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- ALU - operation depends only on the current instruction
--		(decoded in the control unit)
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_arith.all;
use work.p_MR2.all;

entity alu is
	port
	(
		op1, op2: in reg32;
		outalu: out reg32;
		op_alu: in inst_type
	);
end alu;

architecture alu of alu is
	signal menorU, menorS: std_logic;
begin
	menorU <=  '1' when op1 < op2 else '0';
	menorS <=  '1' when IEEE.std_logic_signed."<"(op1, op2) else '0'; -- signed
	outalu <=  op1 - op2
				when  op_alu=SUBU					else
				op1 and op2
				when  op_alu=AAND  or op_alu=ANDI	else
				op1 or  op2
				when  op_alu=OOR	or op_alu=ORI	else
				op1 xor op2
				when  op_alu=XXOR  or op_alu=XORI	else
				to_StdLogicVector(to_bitvector(op1) sll
				CONV_INTEGER(op2(10 downto 6)))
				when  op_alu=SSLL					else
				to_StdLogicVector(to_bitvector(op1) srl
				CONV_INTEGER(op2(10 downto 6)))
				when  op_alu=SSRL					else
				op2(15 downto 0) & x"0000"
				when  op_alu=LUI					else
				(0 => menorU, others => '0')
				when  op_alu=SLTU or op_alu=SLTIU	else	-- signed
				(0 => menorS, others => '0')
				when  op_alu=SLT  or op_alu=SLTI	else	-- unsigned
				-- 22/11/2004 - subtle error correctionwas done for J!
				-- Part of the work for J has been done before, by shifting IR(15 downto 0)
				-- left by two bits before writing data to the IMED register
				op1(31 downto 28) & op2(27 downto 0)
					when  op_alu=J					else
				op1
					when  op_alu=JR	or op_alu=JALR	else
				op1 + op2;
				-- default for ADDU,ADDIU,LBU,LW,SW,SB,BEQ,BGEZ,BLEZ,BNE
end alu;

-------------------------------------------------------------------------
-- Datapath structural description
-------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all; -- needed for comparison instructions SLTxx
use work.p_MR2.all;

entity datapath is
	port
	(
		ck, rst: in std_logic;
		i_address: out reg32;
		instruction: in reg32;
		d_address: out reg32;
		data: inout reg32;
		uins: in microinstruction;
		IR_OUT:	out reg32
	);
end datapath;

architecture datapath of datapath is

	signal incpc, pc, npc, IR,  result, R1, R2, RS, RT, RIN,
			ext16, cte_im, IMED, op1, op2, outalu, RALU, MDR,
			mdr_int, dtpc: reg32 := (others =>  '0');
	signal adD, adS: std_logic_vector(4 downto 0):= (others => '0');
	signal inst_branch, inst_grupo1, inst_grupoI: std_logic;
	signal salta: std_logic:= '0';
	alias ixRS: std_logic_vector(4 downto 0) is IR(25 downto 21);	--  index to Rs --
	alias ixRT: std_logic_vector(4 downto 0) is IR(20 downto 16);	--  index to Rt --

begin

	-- auxiliary signals
	inst_branch <= '1' when uins.i=BEQ or uins.i=BGEZ or uins.i=BLEZ or uins.i=BNE else
				'0';
	inst_grupo1 <= '1' when uins.i=ADDU or uins.i=SUBU or uins.i=AAND or uins.i=OOR or uins.i=XXOR else
				'0';
	inst_grupoI <= '1' when uins.i=ADDIU or uins.i=ANDI or uins.i=ORI or uins.i=XORI else
				'0';

	--==============================================================================
	-- first_stage
	--==============================================================================

	incpc <= pc + 4;
	RNPC: entity work.regnbit generic map(N=>32) port map(ck=>ck, rst=>rst, ce=>uins.CY1, D=>incpc, Q=>npc);
	RIR:  entity work.regnbit generic map(N=>32) port map(ck=>ck, rst=>rst, ce=>uins.CY1, D=>instruction, Q=>IR);
	IR_OUT <= ir;	-- IR is the datapath output signal to carry the instruction
	i_address <= pc;  -- connects PC output to the instruction memory address bus

	--==============================================================================
	-- second stage
	--==============================================================================

	-- signal to be written into the register bank
	RIN <= npc when uins.i=JALR else result;

	-- register bank write address selection
	adD <= 	IR(15 downto 11) when inst_grupo1='1' or uins.i=SLTU or uins.i=SLT or uins.i=JALR else
			IR(20 downto 16); -- inst_grupoI='1' or uins.i=SLTIU or uins.i=SLTI or uins.i=LW or  uins.i=LBU  or uins.i=LUI, or default

	adS <= IR(20 downto 16) when uins.i=SSLL or uins.i=SSRL else -- only for shifts
	       IR(25 downto 21); -- this is the default

	REGS: entity work.reg_bank port map (ck => ck, rst => rst, wreg => uins.wreg, AdRs => adS, AdRt => ir(20 downto 16), adRD => adD, RD => RIN, R1 => R1, R2 => R2);
	-- sign extension
	ext16 <= x"FFFF" & IR(15 downto 0) when IR(15)='1' else x"0000" & IR(15 downto 0);
	-- Immediate constant
	cte_im <= ext16(29 downto 0)  & "00"	when inst_branch='1'	else
			-- branch address adjustment for word frontier
			"0000" & IR(25 downto 0) & "00" when uins.i=J  else
				-- J is word addressed. MSB four bits are defined at the ALU, not here!
			x"0000" & IR(15 downto 0) when uins.i=ANDI or uins.i=ORI or uins.i=XORI else
				-- logic instructions with immediate operand are zero extended
			ext16;
				-- The default case is used by addiu, lbu, lw, sbu and sw instructions
	-- second stage registers
	REG_A:  entity work.regnbit generic map(N=>32) port map(ck=>ck, rst=>rst, ce=>uins.CY2, D=>R1,	    Q=>RS);
	REG_B:  entity work.regnbit generic map(N=>32) port map(ck=>ck, rst=>rst, ce=>uins.CY2, D=>R2,	    Q=>RT);
	REG_IM: entity work.regnbit generic map(N=>32) port map(ck=>ck, rst=>rst, ce=>uins.CY2, D=>cte_im, Q=>IMED);

  --==============================================================================
	-- third stage
	--==============================================================================

	-- select the first ALU operand
	op1 <= pc when inst_branch='1' else	RS;
	-- select the second ALU operand
	op2 <= RT when inst_grupo1='1' or uins.i=SLTU or uins.i=SLT or uins.i=JR else IMED;
	-- ALU instantiation
	inst_alu: entity work.alu port map(op1 => op1, op2 => op2, outalu => outalu, op_alu => uins.i);
	-- ALU registes
	REG_alu: entity work.regnbit generic map(N=>32) port map(ck=>ck, rst=>rst, ce=>uins.wula, D=>outalu, Q=>RALU);
	-- contition to take the branch instructions
	salta <= '1' when ( (RS=RT  and uins.i=BEQ)  or (RS>=0  and uins.i=BGEZ) or
					    (RS <= 0  and uins.i=BLEZ) or (RS/=RT and uins.i=BNE) )  else
			'0';
	result <= MDR when uins.i=LW or uins.i=LBU else RALU;

	--==============================================================================
	-- fourth stage
	--==============================================================================

	d_address <= RALU;
	-- tristate to control memory write
	data <= RT when (uins.ceRW='1' and uins.rw='0') else (others => 'Z');

	-- single byte reading from memory
	mdr_int <= data when uins.i=LW  else x"000000" & data(7 downto 0);
	RMDR: entity work.regnbit generic map(N=>32) port map(ck=>ck, rst=>rst, ce=>uins.wmdr, D=>mdr_int, Q=>MDR);

	--==============================================================================
	-- fifth stage
	--==============================================================================

	dtpc <= result when (inst_branch='1' and salta='1') or uins.i=J or uins.i=JALR or uins.i=JR  else npc;

	--  Data memory starting address: beware of the OFFSET!
	rpc: entity work.regnbit generic map(N=>32, INIT_VALUE=>x"00400000") port map(ck=>ck, rst=>rst, ce=>uins.wpc, D=>dtpc, Q=>pc);

end datapath;

-------------------------------------------------------------------------
--  Control Unit behavioral description
--------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.p_MR2.all;

entity control_unit is
	port
	(
		ck, rst: in std_logic;
		uins: out microinstruction;
		ir: in reg32
	);
end control_unit;

architecture control_unit of control_unit is
	type type_state is (Sidle, Sfetch, Sreg, Salu, Wbk, Sld, Sst, Salta);
	signal em_andamento: std_logic;
	signal EA, PE: type_state;
	signal i: inst_type;
begin
	----------------------------------------------------------------------------------------
	-- BLOCK (1/3) - INSTRUCTION DECODING and ALU operation definition.
	-- This block generates 1 Output Function of the Control Unit
	----------------------------------------------------------------------------------------
	i <=	ADDU  when ir(31 downto 26)="000000" and ir(5 downto 0)="100001" else
			SUBU  when ir(31 downto 26)="000000" and ir(5 downto 0)="100011" else
			AAND  when ir(31 downto 26)="000000" and ir(5 downto 0)="100100" else
			OOR   when ir(31 downto 26)="000000" and ir(5 downto 0)="100101" else
			XXOR  when ir(31 downto 26)="000000" and ir(5 downto 0)="100110" else
			SSLL  when ir(31 downto 21)="00000000000" and ir(5 downto 0)="000000" else
			SSRL  when ir(31 downto 21)="00000000000" and ir(5 downto 0)="000010" else
			ADDIU when ir(31 downto 26)="001001" else
			ANDI  when ir(31 downto 26)="001100" else
			ORI   when ir(31 downto 26)="001101" else
			XORI  when ir(31 downto 26)="001110" else
			LUI   when ir(31 downto 26)="001111" else
			LW    when ir(31 downto 26)="100011" else
			LBU   when ir(31 downto 26)="100100" else
			SW    when ir(31 downto 26)="101011" else
			SB    when ir(31 downto 26)="101000" else
			SLTU  when ir(31 downto 26)="000000" and ir(5 downto 0)="101011" else
			SLT   when ir(31 downto 26)="000000" and ir(5 downto 0)="101010" else
			SLTIU when ir(31 downto 26)="001011" else
			SLTI  when ir(31 downto 26)="001010" else
			BEQ   when ir(31 downto 26)="000100" else
			BGEZ  when ir(31 downto 26)="000001" else
			BLEZ  when ir(31 downto 26)="000110" else
			BNE   when ir(31 downto 26)="000101" else
			J     when ir(31 downto 26)="000010" else
			JALR  when ir(31 downto 26)="000000"  and ir(20 downto 16)="00000" and ir(10 downto 0) = "00000001001" else
			JR    when ir(31 downto 26)="000000" and ir(5 downto 0)="001000" else
			RFE   when ir=x"42000010" else
			ERET  when ir=x"42000018" else
			invalid_instruction; -- IMPORTANT: default condition is invalid instruction;

	assert i /= invalid_instruction
		report "******************* INVALID INSTRUCTION *************"
		severity error;

	uins.i <= i;	-- this instructs the alu to execute its expected operation, if any

	----------------------------------------------------------------------------------------
	-- BLOCK (3/3) - DATAPATH REGISTERS load control signals generation.
	----------------------------------------------------------------------------------------
	uins.CY1  <= '1' when EA=Sfetch else '0';
	uins.CY2  <= '1' when EA=Sreg else '0';
	uins.wula <= '1' when EA=Salu else '0';
	uins.wmdr <= '1' when EA=Sld  else '0';
	uins.wreg <= '1' when EA=Wbk or (EA=salta and i=JALR) else '0';
	uins.rw   <= '0' when EA=Sst else '1';
	uins.ceRW <= '1' when EA=Sld or EA=Sst else '0';
	uins.bw   <= '0' when (EA=Sst and i=SB) else '1';
	uins.wpc  <= '1' when (EA=Wbk or EA=Sst or EA=Salta) else '0';

	---------------------------------------------------------------------------------------------
	-- BLOCK (2/3) - Sequential part of the control unit - two processes implementing the
	-- Control Unit state register and the next-state (combinational) function
	---------------------------------------------------------------------------------------------
	process(rst, ck)
	begin
		if rst='1' then
			EA <= Sidle;
	-- Sidle is the state the machine stays while processor is being reset
		elsif ck'event and ck='1' then
			if EA=Sidle then
				EA <= Sfetch;
			else
				EA <= PE;
			end if;
		end if;
	end process;

	process(EA, i)
		-- NEXT state: depends on the PRESENT state and on the current instruction
	begin
		case EA is
			when Sidle => PE <= Sidle; -- reset being active, the processor do nothing!
			-- first stage:  read the current instruction
			when Sfetch => PE <= Sreg;
			-- second stage: read the register banck and store the mask (when i=stmsk)
			when Sreg => PE <= Salu;
			-- third stage: alu operation
			when Salu  => if i=LW  or i=LBU then
								PE <= Sld;
						elsif i=SW or i=SB then
								PE <= Sst;
						elsif i=J or i=JALR or i=JR or i=BEQ or i=BGEZ or i=BLEZ  or i=BNE then
								PE <= Salta;
						else
								PE <= Wbk;
						end if;
			-- fourth stage: data memory operation
			when Sld  => 	PE <= Wbk;
			-- fifth clock cycle of most instructions  - GO BACK TO FETCH
			when Sst | Salta | Wbk => PE <= Sfetch;
		end case;
	end process;

end control_unit;

entity LI is
	port (
		
		clock_L1, rst: in std_logic;
		ce, rw, bw: in std_logic;
		d_address: in reg32;
		dados: inout reg32;
		halt: out std_logic;

		ce_L12, rw_L12, bw_L12: out std_logic;
		d_address_out_L12: out reg32;
		halt_L12: in std_logic

	);
end entity LI;

architecture behavioral of LI is

	signal hit_L1: std_logic;

begin


end architecture behavioral;

entity LII is
	port (
		
		clock_L2, rst: in std_logic;
		ce_L12, rw_L12, bw_L12: in std_logic;
		d_address_L12: in reg32;
		dados_L12: inout reg32;
		halt_L12: out std_logic;

		clock_L2M: out std_logic;
		ce_L2M, rw_L2M, bw_L2M: out std_logic;
		d_address_out_L2M: out reg32;
		halt_L2M: in std_logic

	);
end entity LII;

architecture behavioral of LII is

	signal hit_L2: std_logic;

begin
	
	clock_L2M <= clockL2_int;
	divisor: process(clock_L2) 
	begin 
		if(rising_edge(clock_L2)) then 
			
			clockL2_int <= not (clock_L2);
		
		end if; 
	end process divisor; 
	
end architecture behavioral;

entity MP is
	port (
		
		clock_L2M, rst: in std_logic;
		ce_L2M, rw_L2M, bw_L2M: in std_logic;
		d_address_L2M: in reg32;
		dados_L2M: inout reg32;
		halt_L2M: out std_logic

		ce_MP, rw_MP, bw_MP: out std_logic;
		d_address_out_MP: out reg32
	);
end entity MP;

architecture behavioral of MP is

begin
	
	divisor: process(clock_L2M) 
	begin 
		if(rising_edge(clock_L2M)) then 

			clockL2M_int <= not(clock_L2M);
		
		end if; 
	end process divisor; 
	
end architecture behavioral;

-------------------------------------------------------------------------
-- Top-level instantiation of the MR2 Datapath and Control Unit
--------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.p_MR2.all;

entity MR2 is
	port
	(
		clock,reset: in std_logic;
		ce: out std_logic_vector(16 downto 0);
		rw, bw: out std_logic;
		i_address, d_address: out reg32;
		instruction: in reg32;
		data: inout reg32;
		intr: in std_logic;
		inta: out std_logic
	);
end MR2;

architecture MR2 of MR2 is
	signal IR: reg32;
	signal uins: microinstruction;
	signal data_address: reg32;
begin

	dp: entity work.datapath port map
	(
		ck => clock,
		rst => reset,
		IR_OUT => IR,
		uins => uins,
		i_address => i_address,
		instruction => instruction,
		d_address => data_address,
		data => data
	);
	ct: entity work.control_unit port map
	(
		ck => clock,
		rst => reset, 
		IR => IR,
		halt => halt,
		uins => uins
	);

	L1: entity work.LI port map (
		
		clock_L1=>clock, rst=>reset,
		ce=>uins.ceRW, rw=>uins.rw, bw=>uins.bw,
		d_address=>data_address, dados=>data,
		halt=>halt,

		ce_L12=>ce_L12, rw_L12=>rw_L12, bw_L12=>bw_L12,
		d_address_out_L12=>d_address_out_L12,
		halt_L12=>halt_L12

	);

	L2: entity work.LII port map (
		
		clock_L2=>clock, rst=>reset,
		ce_L12=>ce_L12, rw_L12=>rw_L12, bw_L12=>bw_L12,
		d_address_L12=>d_address_out_L12, dados_L12=>data,
		halt_L12=>halt_L12,

		clock_L2M=>clock_L2M,
		ce_L2M=>ce_L2M, rw_L2M=>rw_L2M, bw_L2M=>bw_L2M,
		d_address_out_L2M=>d_address_out_L2M,
		halt_L2M=>halt_L2M
	);

	MP: entity work.MP port map (
		
		clock_L2M=>clock_L2M, rst=.reset,
		ce_L2M=>ce_L2M, rw_L2M=>rw_L2M, bw_L2M=>bw_L2M,
		d_address_L2M=>d_address_out_L2M, dados_L2M=>data,
		halt_L2M=>halt_L2M,

		ce_MP=>ce_MP, rw_MP=>rw_MP, bw_MP=>bw_MP,
		d_address_out_MP=>d_address_out_MP
	);

	rw <= rw_MP;
	bw <= bw_MP;

	----------------------------------------------------------------------------------------------------------
	--- Trecho de codigo inserido para habilitar o CE dos periféricos e memória.
	--- 	O ce(0) e da UART
	--- 	O ce(16) e da memória de dados
	--- 	Os demais sao de periféricos de 1 a 15
	--- Alem deste trecho foi inserido a mais na versao gold da MR2:
	---		"APENAS" a codificao da instrucao ERET
	---	Alteracao na entidade com os novos sinais "intr", "inta" e o "ce" de 17 linhas
	----------------------------------------------------------------------------------------------------------
	d_address <= d_address_out_MP;

	ce(0)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE00000" and data_address<x"FFE10000")) else '0';
	ce(1)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE10000" and data_address<x"FFE20000")) else '0';
	ce(2)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE20000" and data_address<x"FFE30000")) else '0';
	ce(3)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE30000" and data_address<x"FFE40000")) else '0';
	ce(4)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE40000" and data_address<x"FFE50000")) else '0';
	ce(5)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE50000" and data_address<x"FFE60000")) else '0';
	ce(6)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE60000" and data_address<x"FFE70000")) else '0';
	ce(7)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE70000" and data_address<x"FFE80000")) else '0';
	ce(8)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE80000" and data_address<x"FFE90000")) else '0';
	ce(9)  <= '1' when (uins.ceRW='1' and (data_address>=x"FFE90000" and data_address<x"FFEA0000")) else '0';
	ce(10) <= '1' when (uins.ceRW='1' and (data_address>=x"FFEA0000" and data_address<x"FFEB0000")) else '0';
	ce(11) <= '1' when (uins.ceRW='1' and (data_address>=x"FFEB0000" and data_address<x"FFEC0000")) else '0';
	ce(12) <= '1' when (uins.ceRW='1' and (data_address>=x"FFEC0000" and data_address<x"FFED0000")) else '0';
	ce(13) <= '1' when (uins.ceRW='1' and (data_address>=x"FFED0000" and data_address<x"FFEE0000")) else '0';
	ce(14) <= '1' when (uins.ceRW='1' and (data_address>=x"FFEE0000" and data_address<x"FFEF0000")) else '0';
	ce(15) <= '1' when (uins.ceRW='1' and (data_address>=x"FFEF0000" and data_address<x"FFF00000")) else '0';
	ce(16) <= '1' when (uins.ceRW='1' and (data_address<x"FFE00000"  or  data_address>=x"FFF00000")) else '0';

end MR2;
